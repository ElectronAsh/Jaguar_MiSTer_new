��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���C	�i��EM'XGi���ozmo��L@��i�ʉ�f�wkmrsuڟ�6A3��ؐ����#�#ߺ��,�^#�+M3��a����?�@���jK�£�_��"kbN�J�/� q�h!�Fm� �,+���)�~��$o����.t�C�Y�C�Q��7�8�p2s�쵿�׎�㏨=����ҵD.����O"�p� @Z�0��ļ"H�H��ӽ���rm�O�L�A��u)���F���'�ý=4��X3�:��
I7�tȱ�%�7���aV��J�)b�piy�gT�f_@�G�rAR��7B���X�Y"^�#�S�Uw�ר`�s�P���U�;e�����Sd�ݾŖi��9)�f97$���t���j���?4�!�7�rM��>����+�>�B y|.iq�L�j�P\� )�w̌���lr�p����fK �p��9-�M,F�ܲҖRb��a/K���R/].��_R�{e����8�?;�9����-�<ꪉA^��1��6�4��p�e歋T-��`����c$ΈR��"�O�y�}����O���%�	���]d��x.Hf��)AǪ��r�ύ����]mF�����<��ֶ�_����E)��q�}��`1�&/g͖��h&I�-E;Ф��'��y��:$���B��{/М*�z$��{�xu��SU���j�����f� ����x��6�b�S{$�#J�Ƅ�WS�&���K�ٻ[\�YB��K��;����s��]1X���>�N�8��� Ry��1�;�� �D��#�����[H���S�Qp�q;�Q�E�D�[����5��m���]�1-����p�o&��)�=�$K�eY��:�#ld=�ށ�^��$������y�\2����i<Yc�L#�a�ߟ��C��#��JqR7�aSp�>�R8AC�/v��ze�<з���P���G�����P�e�Q��+����2�E+�6Ih�Y��Fs`�Yar�*�.��L�bu����>�<@�3t�����L�`�\oq\��I'��	��h��(9#��YOs0�:�u,�k��&q��66d�8�{��?��%���1�c�����fo����O�]�*M�L,�+ѐj�l�i��F=�Heտ3���h2��ߵ���4{}���%\��Li>�sO�1*�{�q�j���)�^ՁV�.kDd,DQ���XN����_hC1���'�(*B�Z&�Fx�YY%S���
MhTL<��a�Z�w]����DmZ���1sYshyM4�;9~Ys�f!�R�1�� ��^�7�R_U���@�5����VXӵ�����Z3�VK�+2E���,� ��ޟ:7����w��7N�U��x�C�zb�$��!M�����ݕ��V��-@�à"�sQ���eTKb�kB����������ⰬH���Y��|�ݹ"p�_k`��G��Bg^��Af��S���o6L�Ǯ��|d�����bW��2�<�kxBvfoA%Q����9���@,FW�$���@�r�0mg�n�>)0wV�	C�96D�<mv��A�-x�N�kW�����[�ٲ�Ei�Cx�5�{hu�Z�@B{L��oB��\�T�+��I'UJ�
J�O����F
��t��ǅ���e��
_��Y'�o-ƆGu� .4B��1�dG�߅�5ZL-{�����D���]=��G��VҖ$d�����<�ŝX�6��Я��Z���C#4W� +|������� �DFaL=��K|L���?��'�~<`�$ �w<����PdR����3'E������0��F�c�9		o�"Iu��'-��L@�<]���`���F��%��&���X���ϗy��0�n���#.���u1�)�+)����tO��˔� �*� �af�ә@�pF��d����*�ڐn� yv+4�D���h�>\���Z��[�5.հ�1Y����7K
pI�ҧ�W8,h�zxN=nds��KG�Ҏ��H���� �	ֆZ4���.=Sīn�o��&$ճ3��_ld���c�h�����I�_Ӳ����~1jS�S@��60��h+�`�X�K$k�m��L��?��P�9^i�J�R�y\m/� �*z9���g}��p����������F�i\��`��gm��z���$��\�	����9���X�/;�;�e�>��������ɑG�� i��p���S�� 